LIBRARY ieee;
use ieee.std_logic_1164.all;
USE IEEE.numeric_std.ALL;
USE IEEE.std_logic_UNSIGNED.ALL;

library work;
use work.trb_net_std.all;
use work.trb_net_components.all;
use work.trb_net16_hub_func.all;
--use work.version.all;

use work.trb_net_gbe_components.all;
use work.trb_net_gbe_protocols.all;

entity gbe_setup is
port(
	CLK                       : in std_logic;
	RESET                     : in std_logic;

	-- interface to regio bus
	BUS_ADDR_IN               : in std_logic_vector(7 downto 0);
	BUS_DATA_IN               : in std_logic_vector(31 downto 0);
	BUS_DATA_OUT              : out std_logic_vector(31 downto 0);
	BUS_WRITE_EN_IN           : in std_logic;
	BUS_READ_EN_IN            : in std_logic;
	BUS_ACK_OUT               : out std_logic;

	-- output to gbe_buf
	GBE_SUBEVENT_ID_OUT       : out std_logic_vector(31 downto 0);
	GBE_SUBEVENT_DEC_OUT      : out std_logic_vector(31 downto 0);
	GBE_QUEUE_DEC_OUT         : out std_logic_vector(31 downto 0);
	GBE_MAX_FRAME_OUT         : out std_logic_vector(15 downto 0);
	GBE_USE_GBE_OUT           : out std_logic;
	GBE_USE_TRBNET_OUT        : out std_logic;
	GBE_USE_MULTIEVENTS_OUT   : out std_logic;
	GBE_READOUT_CTR_OUT       : out std_logic_vector(23 downto 0);
	GBE_READOUT_CTR_VALID_OUT : out std_logic;
	GBE_ALLOW_RX_OUT          : out std_logic;
	GBE_ADDITIONAL_HDR_OUT    : out std_logic;
	GBE_INSERT_TTYPE_OUT      : out std_logic;
	
	MONITOR_RX_BYTES_IN       : in std_logic_vector(31 downto 0);
	MONITOR_RX_FRAMES_IN      : in std_logic_vector(31 downto 0);
	MONITOR_TX_BYTES_IN       : in std_logic_vector(31 downto 0);
	MONITOR_TX_FRAMES_IN      : in std_logic_vector(31 downto 0);
	MONITOR_TX_PACKETS_IN     : in std_logic_vector(31 downto 0);
	MONITOR_DROPPED_IN        : in std_logic_vector(31 downto 0);
	
	MONITOR_SELECT_REC_IN	      : in	std_logic_vector(c_MAX_PROTOCOLS * 32 - 1 downto 0);
	MONITOR_SELECT_REC_BYTES_IN   : in	std_logic_vector(c_MAX_PROTOCOLS * 32 - 1 downto 0);
	MONITOR_SELECT_SENT_BYTES_IN  : in	std_logic_vector(c_MAX_PROTOCOLS * 32 - 1 downto 0);
	MONITOR_SELECT_SENT_IN	      : in	std_logic_vector(c_MAX_PROTOCOLS * 32 - 1 downto 0)
);
end entity;

architecture gbe_setup of gbe_setup is

signal reset_values      : std_logic;
signal subevent_id       : std_logic_vector(31 downto 0);
signal subevent_dec      : std_logic_vector(31 downto 0);
signal queue_dec         : std_logic_vector(31 downto 0);
signal max_frame         : std_logic_vector(15 downto 0);
signal use_gbe           : std_logic;
signal use_trbnet        : std_logic;
signal use_multievents   : std_logic;
signal readout_ctr       : std_logic_vector(23 downto 0);
signal readout_ctr_valid : std_logic;
signal ack               : std_logic;
signal ack_q             : std_logic;
signal data_out          : std_logic_vector(31 downto 0);
signal allow_rx          : std_logic;
signal additional_hdr    : std_logic;
signal insert_ttype      : std_logic;

begin

OUT_PROC : process(CLK)
begin
	if rising_edge(CLK) then
		GBE_SUBEVENT_ID_OUT       <= subevent_id;
		GBE_SUBEVENT_DEC_OUT      <= subevent_dec;
		GBE_QUEUE_DEC_OUT         <= queue_dec;
		GBE_MAX_FRAME_OUT         <= max_frame;
		GBE_USE_GBE_OUT           <= use_gbe;
		GBE_USE_TRBNET_OUT        <= use_trbnet;
		GBE_USE_MULTIEVENTS_OUT   <= use_multievents;
		GBE_READOUT_CTR_OUT       <= readout_ctr;
		GBE_READOUT_CTR_VALID_OUT <= readout_ctr_valid;
		BUS_ACK_OUT               <= ack_q;
		ack_q                     <= ack;
		BUS_DATA_OUT              <= data_out;
		GBE_ALLOW_RX_OUT          <= '1'; --allow_rx;
		GBE_INSERT_TTYPE_OUT      <= insert_ttype;
		GBE_ADDITIONAL_HDR_OUT    <= additional_hdr;
	end if;
end process OUT_PROC;

ACK_PROC : process(CLK)
begin
	if rising_edge(CLK) then
		if (RESET = '1') then
			ack <= '0';
		elsif ((BUS_WRITE_EN_IN = '1') or (BUS_READ_EN_IN = '1')) then
			ack <= '1';
		else
			ack <= '0';
		end if;
	end if;
end process ACK_PROC;

WRITE_PROC : process(CLK)
begin
	if rising_edge(CLK) then
		if ( (RESET = '1') or (reset_values = '1') ) then
			subevent_id       <= x"0000_00cf";
			subevent_dec      <= x"0002_0001";
			queue_dec         <= x"0003_0062";
			max_frame         <= x"0578";
			use_gbe           <= '0';
			use_trbnet        <= '0';
			use_multievents   <= '0';
			reset_values      <= '0';
			readout_ctr       <= x"00_0000";
			readout_ctr_valid <= '0';
			allow_rx          <= '1';
			insert_ttype      <= '0';
			additional_hdr    <= '1';	

		elsif (BUS_WRITE_EN_IN = '1') then
			case BUS_ADDR_IN is

				when x"00" =>
					subevent_id <= BUS_DATA_IN;

				when x"01" =>
					subevent_dec <= BUS_DATA_IN;

				when x"02" =>
					queue_dec <= BUS_DATA_IN;

				when x"04" =>
					max_frame <= BUS_DATA_IN(15 downto 0);
					g_MAX_FRAME_SIZE <= BUS_DATA_IN(15 downto 0);

				when x"05" =>
					if (BUS_DATA_IN = x"0000_0000") then
						use_gbe <= '0';
					else
						use_gbe <= '1';
					end if;

				when x"06" =>
					if (BUS_DATA_IN = x"0000_0000") then
						use_trbnet <= '0';
					else
						use_trbnet <= '1';
					end if;

				when x"07" =>
					if (BUS_DATA_IN = x"0000_0000") then
						use_multievents <= '0';
					else
						use_multievents <= '1';
					end if;

				when x"08" =>
					readout_ctr <= BUS_DATA_IN(23 downto 0);
					readout_ctr_valid <= '1';
					
				when x"09" =>
					allow_rx         <= BUS_DATA_IN(0);
					
				when x"0a" =>
					additional_hdr   <= BUS_DATA_IN(0);
					
				when x"0b" =>
					insert_ttype     <= BUS_DATA_IN(0);

				when x"ff" =>
					if (BUS_DATA_IN = x"ffff_ffff") then
						reset_values <= '1';
					else
						reset_values <= '0';
					end if;

				when others =>
					subevent_id        <= subevent_id;
					subevent_dec       <= subevent_dec;
					queue_dec          <= queue_dec;
					max_frame          <= max_frame;
					use_gbe            <= use_gbe;
					use_trbnet         <= use_trbnet;
					use_multievents    <= use_multievents;
					reset_values       <= reset_values;
					readout_ctr        <= readout_ctr;
					readout_ctr_valid  <= readout_ctr_valid;
					allow_rx           <= allow_rx;
					additional_hdr     <= additional_hdr;
					insert_ttype       <= insert_ttype;
			end case;
		else
			reset_values      <= '0';
			readout_ctr_valid <= '0';
		end if;
	end if;
end process WRITE_PROC;

READ_PROC : process(CLK)
begin
	if rising_edge(CLK) then
		if (RESET = '1') then
			data_out <= (others => '0');
		elsif (BUS_READ_EN_IN = '1') then
			case BUS_ADDR_IN is

				when x"00" =>
					data_out <= subevent_id;

				when x"01" =>
					data_out <= subevent_dec;

				when x"02" =>
					data_out <= queue_dec;

				when x"04" =>
					data_out(15 downto 0) <= max_frame;
					data_out(31 downto 16) <= (others => '0');

				when x"05" =>
					if (use_gbe = '0') then
						data_out <= x"0000_0000";
					else
						data_out <= x"0000_0001";
					end if;

				when x"06" =>
					if (use_trbnet = '0') then
						data_out <= x"0000_0000";
					else
						data_out <= x"0000_0001";
					end if;

				when x"07" =>
					if (use_multievents = '0') then
						data_out <= x"0000_0000";
					else
						data_out <= x"0000_0001";
					end if;
					
				when x"09" =>
					data_out(0) <= allow_rx;
					data_out(31 downto 1) <= (others => '0');
					
				when x"0a" =>
					data_out(0) <= additional_hdr;
					data_out(31 downto 1) <= (others => '0');
					
				when x"0b" =>
					data_out(0) <= insert_ttype;
					data_out(31 downto 1) <= (others => '0');
					
				when x"e0" =>
					data_out <= MONITOR_RX_BYTES_IN;

				when x"e1" =>
					data_out <= MONITOR_RX_FRAMES_IN;

				when x"e2" =>
					data_out <= MONITOR_TX_BYTES_IN;

				when x"e3" =>
					data_out <= MONITOR_TX_FRAMES_IN;

				when x"e4" =>
					data_out <= MONITOR_TX_PACKETS_IN;

				when x"e5" =>
					data_out <= MONITOR_DROPPED_IN;
					
				-- Sctrl
				when x"a0" =>
					data_out <= MONITOR_SELECT_REC_IN(3 * 32 - 1 downto 2 * 32);
				when x"a1" =>
					data_out <= MONITOR_SELECT_REC_BYTES_IN(3 * 32 - 1 downto 2 * 32);
				when x"a2" =>
					data_out <= MONITOR_SELECT_SENT_IN(3 * 32 - 1 downto 2 * 32);
				when x"a3" =>
					data_out <= MONITOR_SELECT_SENT_BYTES_IN(3 * 32 - 1 downto 2 * 32);
					
				-- TrbnetData
				when x"b0" =>
					data_out <= MONITOR_SELECT_REC_IN(4 * 32 - 1 downto 3 * 32);
				when x"b1" =>
					data_out <= MONITOR_SELECT_REC_BYTES_IN(4 * 32 - 1 downto 3 * 32);
				when x"b2" =>
					data_out <= MONITOR_SELECT_SENT_IN(4 * 32 - 1 downto 3 * 32);
				when x"b3" =>
					data_out <= MONITOR_SELECT_SENT_BYTES_IN(4 * 32 - 1 downto 3 * 32);
				
				-- for older network monitors	
				when x"f3" =>
					data_out <= MONITOR_TX_BYTES_IN;
					
				when x"f4" =>
					data_out <= MONITOR_TX_FRAMES_IN;
					
				when others =>
					data_out <= (others => '0');
			end case;
		end if;
	end if;
end process READ_PROC;

end architecture;